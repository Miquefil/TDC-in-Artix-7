
// THIS MODULE HAS BEEN GENERATED WITH THE HELP OF A SCRIPT


module Start_Stop_FlipFlops( 
       input  wire        clk,
       input  wire        iStartEnable,
       input  wire        iStopEnable,
       input  wire        iRst,
      input  wire        [280-1:0] wFirstFF, 
      output wire        [280-1:0] oFFStart, 
      output wire        [280-1:0] oFFStop
); 


(* LOC = "SLICE_X85Y111" *)
      FDCE #(.INIT(1'b0)) Startff0(
          .Q          (oFFStart[0]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[0])
);

(* LOC = "SLICE_X85Y111" *)
      FDCE #(.INIT(1'b0)) Startff1(
          .Q          (oFFStart[1]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[1])
);

(* LOC = "SLICE_X85Y111" *)
      FDCE #(.INIT(1'b0)) Startff2(
          .Q          (oFFStart[2]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[2])
);

(* LOC = "SLICE_X85Y111" *)
      FDCE #(.INIT(1'b0)) Startff3(
          .Q          (oFFStart[3]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[3])
);

(* LOC = "SLICE_X85Y112" *)
      FDCE #(.INIT(1'b0)) Startff4(
          .Q          (oFFStart[4]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[4])
);

(* LOC = "SLICE_X85Y112" *)
      FDCE #(.INIT(1'b0)) Startff5(
          .Q          (oFFStart[5]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[5])
);

(* LOC = "SLICE_X85Y112" *)
      FDCE #(.INIT(1'b0)) Startff6(
          .Q          (oFFStart[6]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[6])
);

(* LOC = "SLICE_X85Y112" *)
      FDCE #(.INIT(1'b0)) Startff7(
          .Q          (oFFStart[7]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[7])
);

(* LOC = "SLICE_X85Y113" *)
      FDCE #(.INIT(1'b0)) Startff8(
          .Q          (oFFStart[8]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[8])
);

(* LOC = "SLICE_X85Y113" *)
      FDCE #(.INIT(1'b0)) Startff9(
          .Q          (oFFStart[9]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[9])
);

(* LOC = "SLICE_X85Y113" *)
      FDCE #(.INIT(1'b0)) Startff10(
          .Q          (oFFStart[10]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[10])
);

(* LOC = "SLICE_X85Y113" *)
      FDCE #(.INIT(1'b0)) Startff11(
          .Q          (oFFStart[11]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[11])
);

(* LOC = "SLICE_X85Y114" *)
      FDCE #(.INIT(1'b0)) Startff12(
          .Q          (oFFStart[12]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[12])
);

(* LOC = "SLICE_X85Y114" *)
      FDCE #(.INIT(1'b0)) Startff13(
          .Q          (oFFStart[13]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[13])
);

(* LOC = "SLICE_X85Y114" *)
      FDCE #(.INIT(1'b0)) Startff14(
          .Q          (oFFStart[14]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[14])
);

(* LOC = "SLICE_X85Y114" *)
      FDCE #(.INIT(1'b0)) Startff15(
          .Q          (oFFStart[15]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[15])
);

(* LOC = "SLICE_X85Y115" *)
      FDCE #(.INIT(1'b0)) Startff16(
          .Q          (oFFStart[16]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[16])
);

(* LOC = "SLICE_X85Y115" *)
      FDCE #(.INIT(1'b0)) Startff17(
          .Q          (oFFStart[17]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[17])
);

(* LOC = "SLICE_X85Y115" *)
      FDCE #(.INIT(1'b0)) Startff18(
          .Q          (oFFStart[18]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[18])
);

(* LOC = "SLICE_X85Y115" *)
      FDCE #(.INIT(1'b0)) Startff19(
          .Q          (oFFStart[19]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[19])
);

(* LOC = "SLICE_X85Y116" *)
      FDCE #(.INIT(1'b0)) Startff20(
          .Q          (oFFStart[20]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[20])
);

(* LOC = "SLICE_X85Y116" *)
      FDCE #(.INIT(1'b0)) Startff21(
          .Q          (oFFStart[21]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[21])
);

(* LOC = "SLICE_X85Y116" *)
      FDCE #(.INIT(1'b0)) Startff22(
          .Q          (oFFStart[22]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[22])
);

(* LOC = "SLICE_X85Y116" *)
      FDCE #(.INIT(1'b0)) Startff23(
          .Q          (oFFStart[23]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[23])
);

(* LOC = "SLICE_X85Y117" *)
      FDCE #(.INIT(1'b0)) Startff24(
          .Q          (oFFStart[24]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[24])
);

(* LOC = "SLICE_X85Y117" *)
      FDCE #(.INIT(1'b0)) Startff25(
          .Q          (oFFStart[25]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[25])
);

(* LOC = "SLICE_X85Y117" *)
      FDCE #(.INIT(1'b0)) Startff26(
          .Q          (oFFStart[26]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[26])
);

(* LOC = "SLICE_X85Y117" *)
      FDCE #(.INIT(1'b0)) Startff27(
          .Q          (oFFStart[27]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[27])
);

(* LOC = "SLICE_X85Y118" *)
      FDCE #(.INIT(1'b0)) Startff28(
          .Q          (oFFStart[28]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[28])
);

(* LOC = "SLICE_X85Y118" *)
      FDCE #(.INIT(1'b0)) Startff29(
          .Q          (oFFStart[29]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[29])
);

(* LOC = "SLICE_X85Y118" *)
      FDCE #(.INIT(1'b0)) Startff30(
          .Q          (oFFStart[30]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[30])
);

(* LOC = "SLICE_X85Y118" *)
      FDCE #(.INIT(1'b0)) Startff31(
          .Q          (oFFStart[31]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[31])
);

(* LOC = "SLICE_X85Y119" *)
      FDCE #(.INIT(1'b0)) Startff32(
          .Q          (oFFStart[32]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[32])
);

(* LOC = "SLICE_X85Y119" *)
      FDCE #(.INIT(1'b0)) Startff33(
          .Q          (oFFStart[33]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[33])
);

(* LOC = "SLICE_X85Y119" *)
      FDCE #(.INIT(1'b0)) Startff34(
          .Q          (oFFStart[34]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[34])
);

(* LOC = "SLICE_X85Y119" *)
      FDCE #(.INIT(1'b0)) Startff35(
          .Q          (oFFStart[35]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[35])
);

(* LOC = "SLICE_X85Y120" *)
      FDCE #(.INIT(1'b0)) Startff36(
          .Q          (oFFStart[36]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[36])
);

(* LOC = "SLICE_X85Y120" *)
      FDCE #(.INIT(1'b0)) Startff37(
          .Q          (oFFStart[37]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[37])
);

(* LOC = "SLICE_X85Y120" *)
      FDCE #(.INIT(1'b0)) Startff38(
          .Q          (oFFStart[38]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[38])
);

(* LOC = "SLICE_X85Y120" *)
      FDCE #(.INIT(1'b0)) Startff39(
          .Q          (oFFStart[39]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[39])
);

(* LOC = "SLICE_X85Y121" *)
      FDCE #(.INIT(1'b0)) Startff40(
          .Q          (oFFStart[40]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[40])
);

(* LOC = "SLICE_X85Y121" *)
      FDCE #(.INIT(1'b0)) Startff41(
          .Q          (oFFStart[41]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[41])
);

(* LOC = "SLICE_X85Y121" *)
      FDCE #(.INIT(1'b0)) Startff42(
          .Q          (oFFStart[42]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[42])
);

(* LOC = "SLICE_X85Y121" *)
      FDCE #(.INIT(1'b0)) Startff43(
          .Q          (oFFStart[43]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[43])
);

(* LOC = "SLICE_X85Y122" *)
      FDCE #(.INIT(1'b0)) Startff44(
          .Q          (oFFStart[44]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[44])
);

(* LOC = "SLICE_X85Y122" *)
      FDCE #(.INIT(1'b0)) Startff45(
          .Q          (oFFStart[45]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[45])
);

(* LOC = "SLICE_X85Y122" *)
      FDCE #(.INIT(1'b0)) Startff46(
          .Q          (oFFStart[46]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[46])
);

(* LOC = "SLICE_X85Y122" *)
      FDCE #(.INIT(1'b0)) Startff47(
          .Q          (oFFStart[47]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[47])
);

(* LOC = "SLICE_X85Y123" *)
      FDCE #(.INIT(1'b0)) Startff48(
          .Q          (oFFStart[48]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[48])
);

(* LOC = "SLICE_X85Y123" *)
      FDCE #(.INIT(1'b0)) Startff49(
          .Q          (oFFStart[49]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[49])
);

(* LOC = "SLICE_X85Y123" *)
      FDCE #(.INIT(1'b0)) Startff50(
          .Q          (oFFStart[50]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[50])
);

(* LOC = "SLICE_X85Y123" *)
      FDCE #(.INIT(1'b0)) Startff51(
          .Q          (oFFStart[51]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[51])
);

(* LOC = "SLICE_X85Y124" *)
      FDCE #(.INIT(1'b0)) Startff52(
          .Q          (oFFStart[52]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[52])
);

(* LOC = "SLICE_X85Y124" *)
      FDCE #(.INIT(1'b0)) Startff53(
          .Q          (oFFStart[53]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[53])
);

(* LOC = "SLICE_X85Y124" *)
      FDCE #(.INIT(1'b0)) Startff54(
          .Q          (oFFStart[54]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[54])
);

(* LOC = "SLICE_X85Y124" *)
      FDCE #(.INIT(1'b0)) Startff55(
          .Q          (oFFStart[55]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[55])
);

(* LOC = "SLICE_X85Y125" *)
      FDCE #(.INIT(1'b0)) Startff56(
          .Q          (oFFStart[56]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[56])
);

(* LOC = "SLICE_X85Y125" *)
      FDCE #(.INIT(1'b0)) Startff57(
          .Q          (oFFStart[57]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[57])
);

(* LOC = "SLICE_X85Y125" *)
      FDCE #(.INIT(1'b0)) Startff58(
          .Q          (oFFStart[58]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[58])
);

(* LOC = "SLICE_X85Y125" *)
      FDCE #(.INIT(1'b0)) Startff59(
          .Q          (oFFStart[59]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[59])
);

(* LOC = "SLICE_X85Y126" *)
      FDCE #(.INIT(1'b0)) Startff60(
          .Q          (oFFStart[60]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[60])
);

(* LOC = "SLICE_X85Y126" *)
      FDCE #(.INIT(1'b0)) Startff61(
          .Q          (oFFStart[61]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[61])
);

(* LOC = "SLICE_X85Y126" *)
      FDCE #(.INIT(1'b0)) Startff62(
          .Q          (oFFStart[62]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[62])
);

(* LOC = "SLICE_X85Y126" *)
      FDCE #(.INIT(1'b0)) Startff63(
          .Q          (oFFStart[63]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[63])
);

(* LOC = "SLICE_X85Y127" *)
      FDCE #(.INIT(1'b0)) Startff64(
          .Q          (oFFStart[64]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[64])
);

(* LOC = "SLICE_X85Y127" *)
      FDCE #(.INIT(1'b0)) Startff65(
          .Q          (oFFStart[65]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[65])
);

(* LOC = "SLICE_X85Y127" *)
      FDCE #(.INIT(1'b0)) Startff66(
          .Q          (oFFStart[66]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[66])
);

(* LOC = "SLICE_X85Y127" *)
      FDCE #(.INIT(1'b0)) Startff67(
          .Q          (oFFStart[67]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[67])
);

(* LOC = "SLICE_X85Y128" *)
      FDCE #(.INIT(1'b0)) Startff68(
          .Q          (oFFStart[68]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[68])
);

(* LOC = "SLICE_X85Y128" *)
      FDCE #(.INIT(1'b0)) Startff69(
          .Q          (oFFStart[69]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[69])
);

(* LOC = "SLICE_X85Y128" *)
      FDCE #(.INIT(1'b0)) Startff70(
          .Q          (oFFStart[70]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[70])
);

(* LOC = "SLICE_X85Y128" *)
      FDCE #(.INIT(1'b0)) Startff71(
          .Q          (oFFStart[71]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[71])
);

(* LOC = "SLICE_X85Y129" *)
      FDCE #(.INIT(1'b0)) Startff72(
          .Q          (oFFStart[72]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[72])
);

(* LOC = "SLICE_X85Y129" *)
      FDCE #(.INIT(1'b0)) Startff73(
          .Q          (oFFStart[73]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[73])
);

(* LOC = "SLICE_X85Y129" *)
      FDCE #(.INIT(1'b0)) Startff74(
          .Q          (oFFStart[74]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[74])
);

(* LOC = "SLICE_X85Y129" *)
      FDCE #(.INIT(1'b0)) Startff75(
          .Q          (oFFStart[75]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[75])
);

(* LOC = "SLICE_X85Y130" *)
      FDCE #(.INIT(1'b0)) Startff76(
          .Q          (oFFStart[76]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[76])
);

(* LOC = "SLICE_X85Y130" *)
      FDCE #(.INIT(1'b0)) Startff77(
          .Q          (oFFStart[77]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[77])
);

(* LOC = "SLICE_X85Y130" *)
      FDCE #(.INIT(1'b0)) Startff78(
          .Q          (oFFStart[78]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[78])
);

(* LOC = "SLICE_X85Y130" *)
      FDCE #(.INIT(1'b0)) Startff79(
          .Q          (oFFStart[79]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[79])
);

(* LOC = "SLICE_X85Y131" *)
      FDCE #(.INIT(1'b0)) Startff80(
          .Q          (oFFStart[80]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[80])
);

(* LOC = "SLICE_X85Y131" *)
      FDCE #(.INIT(1'b0)) Startff81(
          .Q          (oFFStart[81]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[81])
);

(* LOC = "SLICE_X85Y131" *)
      FDCE #(.INIT(1'b0)) Startff82(
          .Q          (oFFStart[82]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[82])
);

(* LOC = "SLICE_X85Y131" *)
      FDCE #(.INIT(1'b0)) Startff83(
          .Q          (oFFStart[83]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[83])
);

(* LOC = "SLICE_X85Y132" *)
      FDCE #(.INIT(1'b0)) Startff84(
          .Q          (oFFStart[84]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[84])
);

(* LOC = "SLICE_X85Y132" *)
      FDCE #(.INIT(1'b0)) Startff85(
          .Q          (oFFStart[85]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[85])
);

(* LOC = "SLICE_X85Y132" *)
      FDCE #(.INIT(1'b0)) Startff86(
          .Q          (oFFStart[86]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[86])
);

(* LOC = "SLICE_X85Y132" *)
      FDCE #(.INIT(1'b0)) Startff87(
          .Q          (oFFStart[87]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[87])
);

(* LOC = "SLICE_X85Y133" *)
      FDCE #(.INIT(1'b0)) Startff88(
          .Q          (oFFStart[88]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[88])
);

(* LOC = "SLICE_X85Y133" *)
      FDCE #(.INIT(1'b0)) Startff89(
          .Q          (oFFStart[89]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[89])
);

(* LOC = "SLICE_X85Y133" *)
      FDCE #(.INIT(1'b0)) Startff90(
          .Q          (oFFStart[90]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[90])
);

(* LOC = "SLICE_X85Y133" *)
      FDCE #(.INIT(1'b0)) Startff91(
          .Q          (oFFStart[91]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[91])
);

(* LOC = "SLICE_X85Y134" *)
      FDCE #(.INIT(1'b0)) Startff92(
          .Q          (oFFStart[92]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[92])
);

(* LOC = "SLICE_X85Y134" *)
      FDCE #(.INIT(1'b0)) Startff93(
          .Q          (oFFStart[93]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[93])
);

(* LOC = "SLICE_X85Y134" *)
      FDCE #(.INIT(1'b0)) Startff94(
          .Q          (oFFStart[94]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[94])
);

(* LOC = "SLICE_X85Y134" *)
      FDCE #(.INIT(1'b0)) Startff95(
          .Q          (oFFStart[95]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[95])
);

(* LOC = "SLICE_X85Y135" *)
      FDCE #(.INIT(1'b0)) Startff96(
          .Q          (oFFStart[96]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[96])
);

(* LOC = "SLICE_X85Y135" *)
      FDCE #(.INIT(1'b0)) Startff97(
          .Q          (oFFStart[97]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[97])
);

(* LOC = "SLICE_X85Y135" *)
      FDCE #(.INIT(1'b0)) Startff98(
          .Q          (oFFStart[98]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[98])
);

(* LOC = "SLICE_X85Y135" *)
      FDCE #(.INIT(1'b0)) Startff99(
          .Q          (oFFStart[99]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[99])
);

(* LOC = "SLICE_X85Y136" *)
      FDCE #(.INIT(1'b0)) Startff100(
          .Q          (oFFStart[100]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[100])
);

(* LOC = "SLICE_X85Y136" *)
      FDCE #(.INIT(1'b0)) Startff101(
          .Q          (oFFStart[101]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[101])
);

(* LOC = "SLICE_X85Y136" *)
      FDCE #(.INIT(1'b0)) Startff102(
          .Q          (oFFStart[102]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[102])
);

(* LOC = "SLICE_X85Y136" *)
      FDCE #(.INIT(1'b0)) Startff103(
          .Q          (oFFStart[103]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[103])
);

(* LOC = "SLICE_X85Y137" *)
      FDCE #(.INIT(1'b0)) Startff104(
          .Q          (oFFStart[104]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[104])
);

(* LOC = "SLICE_X85Y137" *)
      FDCE #(.INIT(1'b0)) Startff105(
          .Q          (oFFStart[105]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[105])
);

(* LOC = "SLICE_X85Y137" *)
      FDCE #(.INIT(1'b0)) Startff106(
          .Q          (oFFStart[106]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[106])
);

(* LOC = "SLICE_X85Y137" *)
      FDCE #(.INIT(1'b0)) Startff107(
          .Q          (oFFStart[107]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[107])
);

(* LOC = "SLICE_X85Y138" *)
      FDCE #(.INIT(1'b0)) Startff108(
          .Q          (oFFStart[108]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[108])
);

(* LOC = "SLICE_X85Y138" *)
      FDCE #(.INIT(1'b0)) Startff109(
          .Q          (oFFStart[109]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[109])
);

(* LOC = "SLICE_X85Y138" *)
      FDCE #(.INIT(1'b0)) Startff110(
          .Q          (oFFStart[110]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[110])
);

(* LOC = "SLICE_X85Y138" *)
      FDCE #(.INIT(1'b0)) Startff111(
          .Q          (oFFStart[111]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[111])
);

(* LOC = "SLICE_X85Y139" *)
      FDCE #(.INIT(1'b0)) Startff112(
          .Q          (oFFStart[112]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[112])
);

(* LOC = "SLICE_X85Y139" *)
      FDCE #(.INIT(1'b0)) Startff113(
          .Q          (oFFStart[113]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[113])
);

(* LOC = "SLICE_X85Y139" *)
      FDCE #(.INIT(1'b0)) Startff114(
          .Q          (oFFStart[114]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[114])
);

(* LOC = "SLICE_X85Y139" *)
      FDCE #(.INIT(1'b0)) Startff115(
          .Q          (oFFStart[115]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[115])
);

(* LOC = "SLICE_X85Y140" *)
      FDCE #(.INIT(1'b0)) Startff116(
          .Q          (oFFStart[116]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[116])
);

(* LOC = "SLICE_X85Y140" *)
      FDCE #(.INIT(1'b0)) Startff117(
          .Q          (oFFStart[117]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[117])
);

(* LOC = "SLICE_X85Y140" *)
      FDCE #(.INIT(1'b0)) Startff118(
          .Q          (oFFStart[118]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[118])
);

(* LOC = "SLICE_X85Y140" *)
      FDCE #(.INIT(1'b0)) Startff119(
          .Q          (oFFStart[119]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[119])
);

(* LOC = "SLICE_X85Y141" *)
      FDCE #(.INIT(1'b0)) Startff120(
          .Q          (oFFStart[120]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[120])
);

(* LOC = "SLICE_X85Y141" *)
      FDCE #(.INIT(1'b0)) Startff121(
          .Q          (oFFStart[121]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[121])
);

(* LOC = "SLICE_X85Y141" *)
      FDCE #(.INIT(1'b0)) Startff122(
          .Q          (oFFStart[122]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[122])
);

(* LOC = "SLICE_X85Y141" *)
      FDCE #(.INIT(1'b0)) Startff123(
          .Q          (oFFStart[123]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[123])
);

(* LOC = "SLICE_X85Y142" *)
      FDCE #(.INIT(1'b0)) Startff124(
          .Q          (oFFStart[124]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[124])
);

(* LOC = "SLICE_X85Y142" *)
      FDCE #(.INIT(1'b0)) Startff125(
          .Q          (oFFStart[125]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[125])
);

(* LOC = "SLICE_X85Y142" *)
      FDCE #(.INIT(1'b0)) Startff126(
          .Q          (oFFStart[126]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[126])
);

(* LOC = "SLICE_X85Y142" *)
      FDCE #(.INIT(1'b0)) Startff127(
          .Q          (oFFStart[127]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[127])
);

(* LOC = "SLICE_X85Y143" *)
      FDCE #(.INIT(1'b0)) Startff128(
          .Q          (oFFStart[128]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[128])
);

(* LOC = "SLICE_X85Y143" *)
      FDCE #(.INIT(1'b0)) Startff129(
          .Q          (oFFStart[129]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[129])
);

(* LOC = "SLICE_X85Y143" *)
      FDCE #(.INIT(1'b0)) Startff130(
          .Q          (oFFStart[130]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[130])
);

(* LOC = "SLICE_X85Y143" *)
      FDCE #(.INIT(1'b0)) Startff131(
          .Q          (oFFStart[131]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[131])
);

(* LOC = "SLICE_X85Y144" *)
      FDCE #(.INIT(1'b0)) Startff132(
          .Q          (oFFStart[132]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[132])
);

(* LOC = "SLICE_X85Y144" *)
      FDCE #(.INIT(1'b0)) Startff133(
          .Q          (oFFStart[133]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[133])
);

(* LOC = "SLICE_X85Y144" *)
      FDCE #(.INIT(1'b0)) Startff134(
          .Q          (oFFStart[134]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[134])
);

(* LOC = "SLICE_X85Y144" *)
      FDCE #(.INIT(1'b0)) Startff135(
          .Q          (oFFStart[135]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[135])
);

(* LOC = "SLICE_X85Y145" *)
      FDCE #(.INIT(1'b0)) Startff136(
          .Q          (oFFStart[136]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[136])
);

(* LOC = "SLICE_X85Y145" *)
      FDCE #(.INIT(1'b0)) Startff137(
          .Q          (oFFStart[137]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[137])
);

(* LOC = "SLICE_X85Y145" *)
      FDCE #(.INIT(1'b0)) Startff138(
          .Q          (oFFStart[138]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[138])
);

(* LOC = "SLICE_X85Y145" *)
      FDCE #(.INIT(1'b0)) Startff139(
          .Q          (oFFStart[139]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[139])
);

(* LOC = "SLICE_X85Y146" *)
      FDCE #(.INIT(1'b0)) Startff140(
          .Q          (oFFStart[140]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[140])
);

(* LOC = "SLICE_X85Y146" *)
      FDCE #(.INIT(1'b0)) Startff141(
          .Q          (oFFStart[141]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[141])
);

(* LOC = "SLICE_X85Y146" *)
      FDCE #(.INIT(1'b0)) Startff142(
          .Q          (oFFStart[142]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[142])
);

(* LOC = "SLICE_X85Y146" *)
      FDCE #(.INIT(1'b0)) Startff143(
          .Q          (oFFStart[143]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[143])
);

(* LOC = "SLICE_X85Y147" *)
      FDCE #(.INIT(1'b0)) Startff144(
          .Q          (oFFStart[144]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[144])
);

(* LOC = "SLICE_X85Y147" *)
      FDCE #(.INIT(1'b0)) Startff145(
          .Q          (oFFStart[145]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[145])
);

(* LOC = "SLICE_X85Y147" *)
      FDCE #(.INIT(1'b0)) Startff146(
          .Q          (oFFStart[146]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[146])
);

(* LOC = "SLICE_X85Y147" *)
      FDCE #(.INIT(1'b0)) Startff147(
          .Q          (oFFStart[147]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[147])
);

(* LOC = "SLICE_X85Y148" *)
      FDCE #(.INIT(1'b0)) Startff148(
          .Q          (oFFStart[148]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[148])
);

(* LOC = "SLICE_X85Y148" *)
      FDCE #(.INIT(1'b0)) Startff149(
          .Q          (oFFStart[149]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[149])
);

(* LOC = "SLICE_X85Y148" *)
      FDCE #(.INIT(1'b0)) Startff150(
          .Q          (oFFStart[150]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[150])
);

(* LOC = "SLICE_X85Y148" *)
      FDCE #(.INIT(1'b0)) Startff151(
          .Q          (oFFStart[151]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[151])
);

(* LOC = "SLICE_X85Y149" *)
      FDCE #(.INIT(1'b0)) Startff152(
          .Q          (oFFStart[152]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[152])
);

(* LOC = "SLICE_X85Y149" *)
      FDCE #(.INIT(1'b0)) Startff153(
          .Q          (oFFStart[153]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[153])
);

(* LOC = "SLICE_X85Y149" *)
      FDCE #(.INIT(1'b0)) Startff154(
          .Q          (oFFStart[154]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[154])
);

(* LOC = "SLICE_X85Y149" *)
      FDCE #(.INIT(1'b0)) Startff155(
          .Q          (oFFStart[155]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[155])
);

(* LOC = "SLICE_X85Y150" *)
      FDCE #(.INIT(1'b0)) Startff156(
          .Q          (oFFStart[156]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[156])
);

(* LOC = "SLICE_X85Y150" *)
      FDCE #(.INIT(1'b0)) Startff157(
          .Q          (oFFStart[157]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[157])
);

(* LOC = "SLICE_X85Y150" *)
      FDCE #(.INIT(1'b0)) Startff158(
          .Q          (oFFStart[158]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[158])
);

(* LOC = "SLICE_X85Y150" *)
      FDCE #(.INIT(1'b0)) Startff159(
          .Q          (oFFStart[159]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[159])
);

(* LOC = "SLICE_X85Y151" *)
      FDCE #(.INIT(1'b0)) Startff160(
          .Q          (oFFStart[160]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[160])
);

(* LOC = "SLICE_X85Y151" *)
      FDCE #(.INIT(1'b0)) Startff161(
          .Q          (oFFStart[161]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[161])
);

(* LOC = "SLICE_X85Y151" *)
      FDCE #(.INIT(1'b0)) Startff162(
          .Q          (oFFStart[162]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[162])
);

(* LOC = "SLICE_X85Y151" *)
      FDCE #(.INIT(1'b0)) Startff163(
          .Q          (oFFStart[163]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[163])
);

(* LOC = "SLICE_X85Y152" *)
      FDCE #(.INIT(1'b0)) Startff164(
          .Q          (oFFStart[164]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[164])
);

(* LOC = "SLICE_X85Y152" *)
      FDCE #(.INIT(1'b0)) Startff165(
          .Q          (oFFStart[165]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[165])
);

(* LOC = "SLICE_X85Y152" *)
      FDCE #(.INIT(1'b0)) Startff166(
          .Q          (oFFStart[166]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[166])
);

(* LOC = "SLICE_X85Y152" *)
      FDCE #(.INIT(1'b0)) Startff167(
          .Q          (oFFStart[167]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[167])
);

(* LOC = "SLICE_X85Y153" *)
      FDCE #(.INIT(1'b0)) Startff168(
          .Q          (oFFStart[168]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[168])
);

(* LOC = "SLICE_X85Y153" *)
      FDCE #(.INIT(1'b0)) Startff169(
          .Q          (oFFStart[169]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[169])
);

(* LOC = "SLICE_X85Y153" *)
      FDCE #(.INIT(1'b0)) Startff170(
          .Q          (oFFStart[170]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[170])
);

(* LOC = "SLICE_X85Y153" *)
      FDCE #(.INIT(1'b0)) Startff171(
          .Q          (oFFStart[171]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[171])
);

(* LOC = "SLICE_X85Y154" *)
      FDCE #(.INIT(1'b0)) Startff172(
          .Q          (oFFStart[172]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[172])
);

(* LOC = "SLICE_X85Y154" *)
      FDCE #(.INIT(1'b0)) Startff173(
          .Q          (oFFStart[173]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[173])
);

(* LOC = "SLICE_X85Y154" *)
      FDCE #(.INIT(1'b0)) Startff174(
          .Q          (oFFStart[174]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[174])
);

(* LOC = "SLICE_X85Y154" *)
      FDCE #(.INIT(1'b0)) Startff175(
          .Q          (oFFStart[175]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[175])
);

(* LOC = "SLICE_X85Y155" *)
      FDCE #(.INIT(1'b0)) Startff176(
          .Q          (oFFStart[176]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[176])
);

(* LOC = "SLICE_X85Y155" *)
      FDCE #(.INIT(1'b0)) Startff177(
          .Q          (oFFStart[177]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[177])
);

(* LOC = "SLICE_X85Y155" *)
      FDCE #(.INIT(1'b0)) Startff178(
          .Q          (oFFStart[178]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[178])
);

(* LOC = "SLICE_X85Y155" *)
      FDCE #(.INIT(1'b0)) Startff179(
          .Q          (oFFStart[179]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[179])
);

(* LOC = "SLICE_X85Y156" *)
      FDCE #(.INIT(1'b0)) Startff180(
          .Q          (oFFStart[180]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[180])
);

(* LOC = "SLICE_X85Y156" *)
      FDCE #(.INIT(1'b0)) Startff181(
          .Q          (oFFStart[181]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[181])
);

(* LOC = "SLICE_X85Y156" *)
      FDCE #(.INIT(1'b0)) Startff182(
          .Q          (oFFStart[182]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[182])
);

(* LOC = "SLICE_X85Y156" *)
      FDCE #(.INIT(1'b0)) Startff183(
          .Q          (oFFStart[183]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[183])
);

(* LOC = "SLICE_X85Y157" *)
      FDCE #(.INIT(1'b0)) Startff184(
          .Q          (oFFStart[184]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[184])
);

(* LOC = "SLICE_X85Y157" *)
      FDCE #(.INIT(1'b0)) Startff185(
          .Q          (oFFStart[185]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[185])
);

(* LOC = "SLICE_X85Y157" *)
      FDCE #(.INIT(1'b0)) Startff186(
          .Q          (oFFStart[186]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[186])
);

(* LOC = "SLICE_X85Y157" *)
      FDCE #(.INIT(1'b0)) Startff187(
          .Q          (oFFStart[187]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[187])
);

(* LOC = "SLICE_X85Y158" *)
      FDCE #(.INIT(1'b0)) Startff188(
          .Q          (oFFStart[188]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[188])
);

(* LOC = "SLICE_X85Y158" *)
      FDCE #(.INIT(1'b0)) Startff189(
          .Q          (oFFStart[189]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[189])
);

(* LOC = "SLICE_X85Y158" *)
      FDCE #(.INIT(1'b0)) Startff190(
          .Q          (oFFStart[190]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[190])
);

(* LOC = "SLICE_X85Y158" *)
      FDCE #(.INIT(1'b0)) Startff191(
          .Q          (oFFStart[191]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[191])
);

(* LOC = "SLICE_X85Y159" *)
      FDCE #(.INIT(1'b0)) Startff192(
          .Q          (oFFStart[192]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[192])
);

(* LOC = "SLICE_X85Y159" *)
      FDCE #(.INIT(1'b0)) Startff193(
          .Q          (oFFStart[193]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[193])
);

(* LOC = "SLICE_X85Y159" *)
      FDCE #(.INIT(1'b0)) Startff194(
          .Q          (oFFStart[194]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[194])
);

(* LOC = "SLICE_X85Y159" *)
      FDCE #(.INIT(1'b0)) Startff195(
          .Q          (oFFStart[195]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[195])
);

(* LOC = "SLICE_X85Y160" *)
      FDCE #(.INIT(1'b0)) Startff196(
          .Q          (oFFStart[196]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[196])
);

(* LOC = "SLICE_X85Y160" *)
      FDCE #(.INIT(1'b0)) Startff197(
          .Q          (oFFStart[197]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[197])
);

(* LOC = "SLICE_X85Y160" *)
      FDCE #(.INIT(1'b0)) Startff198(
          .Q          (oFFStart[198]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[198])
);

(* LOC = "SLICE_X85Y160" *)
      FDCE #(.INIT(1'b0)) Startff199(
          .Q          (oFFStart[199]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[199])
);

(* LOC = "SLICE_X85Y161" *)
      FDCE #(.INIT(1'b0)) Startff200(
          .Q          (oFFStart[200]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[200])
);

(* LOC = "SLICE_X85Y161" *)
      FDCE #(.INIT(1'b0)) Startff201(
          .Q          (oFFStart[201]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[201])
);

(* LOC = "SLICE_X85Y161" *)
      FDCE #(.INIT(1'b0)) Startff202(
          .Q          (oFFStart[202]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[202])
);

(* LOC = "SLICE_X85Y161" *)
      FDCE #(.INIT(1'b0)) Startff203(
          .Q          (oFFStart[203]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[203])
);

(* LOC = "SLICE_X85Y162" *)
      FDCE #(.INIT(1'b0)) Startff204(
          .Q          (oFFStart[204]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[204])
);

(* LOC = "SLICE_X85Y162" *)
      FDCE #(.INIT(1'b0)) Startff205(
          .Q          (oFFStart[205]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[205])
);

(* LOC = "SLICE_X85Y162" *)
      FDCE #(.INIT(1'b0)) Startff206(
          .Q          (oFFStart[206]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[206])
);

(* LOC = "SLICE_X85Y162" *)
      FDCE #(.INIT(1'b0)) Startff207(
          .Q          (oFFStart[207]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[207])
);

(* LOC = "SLICE_X85Y163" *)
      FDCE #(.INIT(1'b0)) Startff208(
          .Q          (oFFStart[208]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[208])
);

(* LOC = "SLICE_X85Y163" *)
      FDCE #(.INIT(1'b0)) Startff209(
          .Q          (oFFStart[209]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[209])
);

(* LOC = "SLICE_X85Y163" *)
      FDCE #(.INIT(1'b0)) Startff210(
          .Q          (oFFStart[210]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[210])
);

(* LOC = "SLICE_X85Y163" *)
      FDCE #(.INIT(1'b0)) Startff211(
          .Q          (oFFStart[211]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[211])
);

(* LOC = "SLICE_X85Y164" *)
      FDCE #(.INIT(1'b0)) Startff212(
          .Q          (oFFStart[212]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[212])
);

(* LOC = "SLICE_X85Y164" *)
      FDCE #(.INIT(1'b0)) Startff213(
          .Q          (oFFStart[213]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[213])
);

(* LOC = "SLICE_X85Y164" *)
      FDCE #(.INIT(1'b0)) Startff214(
          .Q          (oFFStart[214]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[214])
);

(* LOC = "SLICE_X85Y164" *)
      FDCE #(.INIT(1'b0)) Startff215(
          .Q          (oFFStart[215]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[215])
);

(* LOC = "SLICE_X85Y165" *)
      FDCE #(.INIT(1'b0)) Startff216(
          .Q          (oFFStart[216]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[216])
);

(* LOC = "SLICE_X85Y165" *)
      FDCE #(.INIT(1'b0)) Startff217(
          .Q          (oFFStart[217]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[217])
);

(* LOC = "SLICE_X85Y165" *)
      FDCE #(.INIT(1'b0)) Startff218(
          .Q          (oFFStart[218]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[218])
);

(* LOC = "SLICE_X85Y165" *)
      FDCE #(.INIT(1'b0)) Startff219(
          .Q          (oFFStart[219]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[219])
);

(* LOC = "SLICE_X85Y166" *)
      FDCE #(.INIT(1'b0)) Startff220(
          .Q          (oFFStart[220]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[220])
);

(* LOC = "SLICE_X85Y166" *)
      FDCE #(.INIT(1'b0)) Startff221(
          .Q          (oFFStart[221]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[221])
);

(* LOC = "SLICE_X85Y166" *)
      FDCE #(.INIT(1'b0)) Startff222(
          .Q          (oFFStart[222]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[222])
);

(* LOC = "SLICE_X85Y166" *)
      FDCE #(.INIT(1'b0)) Startff223(
          .Q          (oFFStart[223]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[223])
);

(* LOC = "SLICE_X85Y167" *)
      FDCE #(.INIT(1'b0)) Startff224(
          .Q          (oFFStart[224]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[224])
);

(* LOC = "SLICE_X85Y167" *)
      FDCE #(.INIT(1'b0)) Startff225(
          .Q          (oFFStart[225]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[225])
);

(* LOC = "SLICE_X85Y167" *)
      FDCE #(.INIT(1'b0)) Startff226(
          .Q          (oFFStart[226]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[226])
);

(* LOC = "SLICE_X85Y167" *)
      FDCE #(.INIT(1'b0)) Startff227(
          .Q          (oFFStart[227]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[227])
);

(* LOC = "SLICE_X85Y168" *)
      FDCE #(.INIT(1'b0)) Startff228(
          .Q          (oFFStart[228]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[228])
);

(* LOC = "SLICE_X85Y168" *)
      FDCE #(.INIT(1'b0)) Startff229(
          .Q          (oFFStart[229]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[229])
);

(* LOC = "SLICE_X85Y168" *)
      FDCE #(.INIT(1'b0)) Startff230(
          .Q          (oFFStart[230]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[230])
);

(* LOC = "SLICE_X85Y168" *)
      FDCE #(.INIT(1'b0)) Startff231(
          .Q          (oFFStart[231]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[231])
);

(* LOC = "SLICE_X85Y169" *)
      FDCE #(.INIT(1'b0)) Startff232(
          .Q          (oFFStart[232]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[232])
);

(* LOC = "SLICE_X85Y169" *)
      FDCE #(.INIT(1'b0)) Startff233(
          .Q          (oFFStart[233]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[233])
);

(* LOC = "SLICE_X85Y169" *)
      FDCE #(.INIT(1'b0)) Startff234(
          .Q          (oFFStart[234]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[234])
);

(* LOC = "SLICE_X85Y169" *)
      FDCE #(.INIT(1'b0)) Startff235(
          .Q          (oFFStart[235]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[235])
);

(* LOC = "SLICE_X85Y170" *)
      FDCE #(.INIT(1'b0)) Startff236(
          .Q          (oFFStart[236]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[236])
);

(* LOC = "SLICE_X85Y170" *)
      FDCE #(.INIT(1'b0)) Startff237(
          .Q          (oFFStart[237]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[237])
);

(* LOC = "SLICE_X85Y170" *)
      FDCE #(.INIT(1'b0)) Startff238(
          .Q          (oFFStart[238]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[238])
);

(* LOC = "SLICE_X85Y170" *)
      FDCE #(.INIT(1'b0)) Startff239(
          .Q          (oFFStart[239]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[239])
);

(* LOC = "SLICE_X85Y171" *)
      FDCE #(.INIT(1'b0)) Startff240(
          .Q          (oFFStart[240]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[240])
);

(* LOC = "SLICE_X85Y171" *)
      FDCE #(.INIT(1'b0)) Startff241(
          .Q          (oFFStart[241]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[241])
);

(* LOC = "SLICE_X85Y171" *)
      FDCE #(.INIT(1'b0)) Startff242(
          .Q          (oFFStart[242]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[242])
);

(* LOC = "SLICE_X85Y171" *)
      FDCE #(.INIT(1'b0)) Startff243(
          .Q          (oFFStart[243]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[243])
);

(* LOC = "SLICE_X85Y172" *)
      FDCE #(.INIT(1'b0)) Startff244(
          .Q          (oFFStart[244]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[244])
);

(* LOC = "SLICE_X85Y172" *)
      FDCE #(.INIT(1'b0)) Startff245(
          .Q          (oFFStart[245]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[245])
);

(* LOC = "SLICE_X85Y172" *)
      FDCE #(.INIT(1'b0)) Startff246(
          .Q          (oFFStart[246]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[246])
);

(* LOC = "SLICE_X85Y172" *)
      FDCE #(.INIT(1'b0)) Startff247(
          .Q          (oFFStart[247]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[247])
);

(* LOC = "SLICE_X85Y173" *)
      FDCE #(.INIT(1'b0)) Startff248(
          .Q          (oFFStart[248]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[248])
);

(* LOC = "SLICE_X85Y173" *)
      FDCE #(.INIT(1'b0)) Startff249(
          .Q          (oFFStart[249]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[249])
);

(* LOC = "SLICE_X85Y173" *)
      FDCE #(.INIT(1'b0)) Startff250(
          .Q          (oFFStart[250]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[250])
);

(* LOC = "SLICE_X85Y173" *)
      FDCE #(.INIT(1'b0)) Startff251(
          .Q          (oFFStart[251]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[251])
);

(* LOC = "SLICE_X85Y174" *)
      FDCE #(.INIT(1'b0)) Startff252(
          .Q          (oFFStart[252]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[252])
);

(* LOC = "SLICE_X85Y174" *)
      FDCE #(.INIT(1'b0)) Startff253(
          .Q          (oFFStart[253]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[253])
);

(* LOC = "SLICE_X85Y174" *)
      FDCE #(.INIT(1'b0)) Startff254(
          .Q          (oFFStart[254]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[254])
);

(* LOC = "SLICE_X85Y174" *)
      FDCE #(.INIT(1'b0)) Startff255(
          .Q          (oFFStart[255]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[255])
);

(* LOC = "SLICE_X85Y175" *)
      FDCE #(.INIT(1'b0)) Startff256(
          .Q          (oFFStart[256]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[256])
);

(* LOC = "SLICE_X85Y175" *)
      FDCE #(.INIT(1'b0)) Startff257(
          .Q          (oFFStart[257]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[257])
);

(* LOC = "SLICE_X85Y175" *)
      FDCE #(.INIT(1'b0)) Startff258(
          .Q          (oFFStart[258]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[258])
);

(* LOC = "SLICE_X85Y175" *)
      FDCE #(.INIT(1'b0)) Startff259(
          .Q          (oFFStart[259]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[259])
);

(* LOC = "SLICE_X85Y176" *)
      FDCE #(.INIT(1'b0)) Startff260(
          .Q          (oFFStart[260]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[260])
);

(* LOC = "SLICE_X85Y176" *)
      FDCE #(.INIT(1'b0)) Startff261(
          .Q          (oFFStart[261]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[261])
);

(* LOC = "SLICE_X85Y176" *)
      FDCE #(.INIT(1'b0)) Startff262(
          .Q          (oFFStart[262]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[262])
);

(* LOC = "SLICE_X85Y176" *)
      FDCE #(.INIT(1'b0)) Startff263(
          .Q          (oFFStart[263]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[263])
);

(* LOC = "SLICE_X85Y177" *)
      FDCE #(.INIT(1'b0)) Startff264(
          .Q          (oFFStart[264]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[264])
);

(* LOC = "SLICE_X85Y177" *)
      FDCE #(.INIT(1'b0)) Startff265(
          .Q          (oFFStart[265]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[265])
);

(* LOC = "SLICE_X85Y177" *)
      FDCE #(.INIT(1'b0)) Startff266(
          .Q          (oFFStart[266]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[266])
);

(* LOC = "SLICE_X85Y177" *)
      FDCE #(.INIT(1'b0)) Startff267(
          .Q          (oFFStart[267]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[267])
);

(* LOC = "SLICE_X85Y178" *)
      FDCE #(.INIT(1'b0)) Startff268(
          .Q          (oFFStart[268]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[268])
);

(* LOC = "SLICE_X85Y178" *)
      FDCE #(.INIT(1'b0)) Startff269(
          .Q          (oFFStart[269]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[269])
);

(* LOC = "SLICE_X85Y178" *)
      FDCE #(.INIT(1'b0)) Startff270(
          .Q          (oFFStart[270]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[270])
);

(* LOC = "SLICE_X85Y178" *)
      FDCE #(.INIT(1'b0)) Startff271(
          .Q          (oFFStart[271]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[271])
);

(* LOC = "SLICE_X85Y179" *)
      FDCE #(.INIT(1'b0)) Startff272(
          .Q          (oFFStart[272]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[272])
);

(* LOC = "SLICE_X85Y179" *)
      FDCE #(.INIT(1'b0)) Startff273(
          .Q          (oFFStart[273]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[273])
);

(* LOC = "SLICE_X85Y179" *)
      FDCE #(.INIT(1'b0)) Startff274(
          .Q          (oFFStart[274]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[274])
);

(* LOC = "SLICE_X85Y179" *)
      FDCE #(.INIT(1'b0)) Startff275(
          .Q          (oFFStart[275]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[275])
);

(* LOC = "SLICE_X85Y180" *)
      FDCE #(.INIT(1'b0)) Startff276(
          .Q          (oFFStart[276]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[276])
);

(* LOC = "SLICE_X85Y180" *)
      FDCE #(.INIT(1'b0)) Startff277(
          .Q          (oFFStart[277]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[277])
);

(* LOC = "SLICE_X85Y180" *)
      FDCE #(.INIT(1'b0)) Startff278(
          .Q          (oFFStart[278]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[278])
);

(* LOC = "SLICE_X85Y180" *)
      FDCE #(.INIT(1'b0)) Startff279(
          .Q          (oFFStart[279]),
          .C          (clk),
          .CE         (iStartEnable),
          .CLR        (iRst),
          .D          (wFirstFF[279])
);

(* LOC = "SLICE_X87Y111" *)
      FDCE #(.INIT(1'b0)) Stopff0(
          .Q          (oFFStop[0]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[0])
);

(* LOC = "SLICE_X87Y111" *)
      FDCE #(.INIT(1'b0)) Stopff1(
          .Q          (oFFStop[1]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[1])
);

(* LOC = "SLICE_X87Y111" *)
      FDCE #(.INIT(1'b0)) Stopff2(
          .Q          (oFFStop[2]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[2])
);

(* LOC = "SLICE_X87Y111" *)
      FDCE #(.INIT(1'b0)) Stopff3(
          .Q          (oFFStop[3]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[3])
);

(* LOC = "SLICE_X87Y112" *)
      FDCE #(.INIT(1'b0)) Stopff4(
          .Q          (oFFStop[4]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[4])
);

(* LOC = "SLICE_X87Y112" *)
      FDCE #(.INIT(1'b0)) Stopff5(
          .Q          (oFFStop[5]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[5])
);

(* LOC = "SLICE_X87Y112" *)
      FDCE #(.INIT(1'b0)) Stopff6(
          .Q          (oFFStop[6]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[6])
);

(* LOC = "SLICE_X87Y112" *)
      FDCE #(.INIT(1'b0)) Stopff7(
          .Q          (oFFStop[7]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[7])
);

(* LOC = "SLICE_X87Y113" *)
      FDCE #(.INIT(1'b0)) Stopff8(
          .Q          (oFFStop[8]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[8])
);

(* LOC = "SLICE_X87Y113" *)
      FDCE #(.INIT(1'b0)) Stopff9(
          .Q          (oFFStop[9]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[9])
);

(* LOC = "SLICE_X87Y113" *)
      FDCE #(.INIT(1'b0)) Stopff10(
          .Q          (oFFStop[10]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[10])
);

(* LOC = "SLICE_X87Y113" *)
      FDCE #(.INIT(1'b0)) Stopff11(
          .Q          (oFFStop[11]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[11])
);

(* LOC = "SLICE_X87Y114" *)
      FDCE #(.INIT(1'b0)) Stopff12(
          .Q          (oFFStop[12]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[12])
);

(* LOC = "SLICE_X87Y114" *)
      FDCE #(.INIT(1'b0)) Stopff13(
          .Q          (oFFStop[13]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[13])
);

(* LOC = "SLICE_X87Y114" *)
      FDCE #(.INIT(1'b0)) Stopff14(
          .Q          (oFFStop[14]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[14])
);

(* LOC = "SLICE_X87Y114" *)
      FDCE #(.INIT(1'b0)) Stopff15(
          .Q          (oFFStop[15]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[15])
);

(* LOC = "SLICE_X87Y115" *)
      FDCE #(.INIT(1'b0)) Stopff16(
          .Q          (oFFStop[16]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[16])
);

(* LOC = "SLICE_X87Y115" *)
      FDCE #(.INIT(1'b0)) Stopff17(
          .Q          (oFFStop[17]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[17])
);

(* LOC = "SLICE_X87Y115" *)
      FDCE #(.INIT(1'b0)) Stopff18(
          .Q          (oFFStop[18]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[18])
);

(* LOC = "SLICE_X87Y115" *)
      FDCE #(.INIT(1'b0)) Stopff19(
          .Q          (oFFStop[19]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[19])
);

(* LOC = "SLICE_X87Y116" *)
      FDCE #(.INIT(1'b0)) Stopff20(
          .Q          (oFFStop[20]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[20])
);

(* LOC = "SLICE_X87Y116" *)
      FDCE #(.INIT(1'b0)) Stopff21(
          .Q          (oFFStop[21]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[21])
);

(* LOC = "SLICE_X87Y116" *)
      FDCE #(.INIT(1'b0)) Stopff22(
          .Q          (oFFStop[22]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[22])
);

(* LOC = "SLICE_X87Y116" *)
      FDCE #(.INIT(1'b0)) Stopff23(
          .Q          (oFFStop[23]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[23])
);

(* LOC = "SLICE_X87Y117" *)
      FDCE #(.INIT(1'b0)) Stopff24(
          .Q          (oFFStop[24]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[24])
);

(* LOC = "SLICE_X87Y117" *)
      FDCE #(.INIT(1'b0)) Stopff25(
          .Q          (oFFStop[25]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[25])
);

(* LOC = "SLICE_X87Y117" *)
      FDCE #(.INIT(1'b0)) Stopff26(
          .Q          (oFFStop[26]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[26])
);

(* LOC = "SLICE_X87Y117" *)
      FDCE #(.INIT(1'b0)) Stopff27(
          .Q          (oFFStop[27]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[27])
);

(* LOC = "SLICE_X87Y118" *)
      FDCE #(.INIT(1'b0)) Stopff28(
          .Q          (oFFStop[28]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[28])
);

(* LOC = "SLICE_X87Y118" *)
      FDCE #(.INIT(1'b0)) Stopff29(
          .Q          (oFFStop[29]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[29])
);

(* LOC = "SLICE_X87Y118" *)
      FDCE #(.INIT(1'b0)) Stopff30(
          .Q          (oFFStop[30]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[30])
);

(* LOC = "SLICE_X87Y118" *)
      FDCE #(.INIT(1'b0)) Stopff31(
          .Q          (oFFStop[31]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[31])
);

(* LOC = "SLICE_X87Y119" *)
      FDCE #(.INIT(1'b0)) Stopff32(
          .Q          (oFFStop[32]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[32])
);

(* LOC = "SLICE_X87Y119" *)
      FDCE #(.INIT(1'b0)) Stopff33(
          .Q          (oFFStop[33]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[33])
);

(* LOC = "SLICE_X87Y119" *)
      FDCE #(.INIT(1'b0)) Stopff34(
          .Q          (oFFStop[34]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[34])
);

(* LOC = "SLICE_X87Y119" *)
      FDCE #(.INIT(1'b0)) Stopff35(
          .Q          (oFFStop[35]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[35])
);

(* LOC = "SLICE_X87Y120" *)
      FDCE #(.INIT(1'b0)) Stopff36(
          .Q          (oFFStop[36]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[36])
);

(* LOC = "SLICE_X87Y120" *)
      FDCE #(.INIT(1'b0)) Stopff37(
          .Q          (oFFStop[37]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[37])
);

(* LOC = "SLICE_X87Y120" *)
      FDCE #(.INIT(1'b0)) Stopff38(
          .Q          (oFFStop[38]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[38])
);

(* LOC = "SLICE_X87Y120" *)
      FDCE #(.INIT(1'b0)) Stopff39(
          .Q          (oFFStop[39]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[39])
);

(* LOC = "SLICE_X87Y121" *)
      FDCE #(.INIT(1'b0)) Stopff40(
          .Q          (oFFStop[40]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[40])
);

(* LOC = "SLICE_X87Y121" *)
      FDCE #(.INIT(1'b0)) Stopff41(
          .Q          (oFFStop[41]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[41])
);

(* LOC = "SLICE_X87Y121" *)
      FDCE #(.INIT(1'b0)) Stopff42(
          .Q          (oFFStop[42]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[42])
);

(* LOC = "SLICE_X87Y121" *)
      FDCE #(.INIT(1'b0)) Stopff43(
          .Q          (oFFStop[43]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[43])
);

(* LOC = "SLICE_X87Y122" *)
      FDCE #(.INIT(1'b0)) Stopff44(
          .Q          (oFFStop[44]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[44])
);

(* LOC = "SLICE_X87Y122" *)
      FDCE #(.INIT(1'b0)) Stopff45(
          .Q          (oFFStop[45]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[45])
);

(* LOC = "SLICE_X87Y122" *)
      FDCE #(.INIT(1'b0)) Stopff46(
          .Q          (oFFStop[46]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[46])
);

(* LOC = "SLICE_X87Y122" *)
      FDCE #(.INIT(1'b0)) Stopff47(
          .Q          (oFFStop[47]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[47])
);

(* LOC = "SLICE_X87Y123" *)
      FDCE #(.INIT(1'b0)) Stopff48(
          .Q          (oFFStop[48]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[48])
);

(* LOC = "SLICE_X87Y123" *)
      FDCE #(.INIT(1'b0)) Stopff49(
          .Q          (oFFStop[49]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[49])
);

(* LOC = "SLICE_X87Y123" *)
      FDCE #(.INIT(1'b0)) Stopff50(
          .Q          (oFFStop[50]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[50])
);

(* LOC = "SLICE_X87Y123" *)
      FDCE #(.INIT(1'b0)) Stopff51(
          .Q          (oFFStop[51]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[51])
);

(* LOC = "SLICE_X87Y124" *)
      FDCE #(.INIT(1'b0)) Stopff52(
          .Q          (oFFStop[52]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[52])
);

(* LOC = "SLICE_X87Y124" *)
      FDCE #(.INIT(1'b0)) Stopff53(
          .Q          (oFFStop[53]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[53])
);

(* LOC = "SLICE_X87Y124" *)
      FDCE #(.INIT(1'b0)) Stopff54(
          .Q          (oFFStop[54]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[54])
);

(* LOC = "SLICE_X87Y124" *)
      FDCE #(.INIT(1'b0)) Stopff55(
          .Q          (oFFStop[55]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[55])
);

(* LOC = "SLICE_X87Y125" *)
      FDCE #(.INIT(1'b0)) Stopff56(
          .Q          (oFFStop[56]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[56])
);

(* LOC = "SLICE_X87Y125" *)
      FDCE #(.INIT(1'b0)) Stopff57(
          .Q          (oFFStop[57]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[57])
);

(* LOC = "SLICE_X87Y125" *)
      FDCE #(.INIT(1'b0)) Stopff58(
          .Q          (oFFStop[58]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[58])
);

(* LOC = "SLICE_X87Y125" *)
      FDCE #(.INIT(1'b0)) Stopff59(
          .Q          (oFFStop[59]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[59])
);

(* LOC = "SLICE_X87Y126" *)
      FDCE #(.INIT(1'b0)) Stopff60(
          .Q          (oFFStop[60]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[60])
);

(* LOC = "SLICE_X87Y126" *)
      FDCE #(.INIT(1'b0)) Stopff61(
          .Q          (oFFStop[61]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[61])
);

(* LOC = "SLICE_X87Y126" *)
      FDCE #(.INIT(1'b0)) Stopff62(
          .Q          (oFFStop[62]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[62])
);

(* LOC = "SLICE_X87Y126" *)
      FDCE #(.INIT(1'b0)) Stopff63(
          .Q          (oFFStop[63]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[63])
);

(* LOC = "SLICE_X87Y127" *)
      FDCE #(.INIT(1'b0)) Stopff64(
          .Q          (oFFStop[64]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[64])
);

(* LOC = "SLICE_X87Y127" *)
      FDCE #(.INIT(1'b0)) Stopff65(
          .Q          (oFFStop[65]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[65])
);

(* LOC = "SLICE_X87Y127" *)
      FDCE #(.INIT(1'b0)) Stopff66(
          .Q          (oFFStop[66]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[66])
);

(* LOC = "SLICE_X87Y127" *)
      FDCE #(.INIT(1'b0)) Stopff67(
          .Q          (oFFStop[67]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[67])
);

(* LOC = "SLICE_X87Y128" *)
      FDCE #(.INIT(1'b0)) Stopff68(
          .Q          (oFFStop[68]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[68])
);

(* LOC = "SLICE_X87Y128" *)
      FDCE #(.INIT(1'b0)) Stopff69(
          .Q          (oFFStop[69]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[69])
);

(* LOC = "SLICE_X87Y128" *)
      FDCE #(.INIT(1'b0)) Stopff70(
          .Q          (oFFStop[70]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[70])
);

(* LOC = "SLICE_X87Y128" *)
      FDCE #(.INIT(1'b0)) Stopff71(
          .Q          (oFFStop[71]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[71])
);

(* LOC = "SLICE_X87Y129" *)
      FDCE #(.INIT(1'b0)) Stopff72(
          .Q          (oFFStop[72]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[72])
);

(* LOC = "SLICE_X87Y129" *)
      FDCE #(.INIT(1'b0)) Stopff73(
          .Q          (oFFStop[73]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[73])
);

(* LOC = "SLICE_X87Y129" *)
      FDCE #(.INIT(1'b0)) Stopff74(
          .Q          (oFFStop[74]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[74])
);

(* LOC = "SLICE_X87Y129" *)
      FDCE #(.INIT(1'b0)) Stopff75(
          .Q          (oFFStop[75]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[75])
);

(* LOC = "SLICE_X87Y130" *)
      FDCE #(.INIT(1'b0)) Stopff76(
          .Q          (oFFStop[76]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[76])
);

(* LOC = "SLICE_X87Y130" *)
      FDCE #(.INIT(1'b0)) Stopff77(
          .Q          (oFFStop[77]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[77])
);

(* LOC = "SLICE_X87Y130" *)
      FDCE #(.INIT(1'b0)) Stopff78(
          .Q          (oFFStop[78]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[78])
);

(* LOC = "SLICE_X87Y130" *)
      FDCE #(.INIT(1'b0)) Stopff79(
          .Q          (oFFStop[79]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[79])
);

(* LOC = "SLICE_X87Y131" *)
      FDCE #(.INIT(1'b0)) Stopff80(
          .Q          (oFFStop[80]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[80])
);

(* LOC = "SLICE_X87Y131" *)
      FDCE #(.INIT(1'b0)) Stopff81(
          .Q          (oFFStop[81]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[81])
);

(* LOC = "SLICE_X87Y131" *)
      FDCE #(.INIT(1'b0)) Stopff82(
          .Q          (oFFStop[82]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[82])
);

(* LOC = "SLICE_X87Y131" *)
      FDCE #(.INIT(1'b0)) Stopff83(
          .Q          (oFFStop[83]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[83])
);

(* LOC = "SLICE_X87Y132" *)
      FDCE #(.INIT(1'b0)) Stopff84(
          .Q          (oFFStop[84]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[84])
);

(* LOC = "SLICE_X87Y132" *)
      FDCE #(.INIT(1'b0)) Stopff85(
          .Q          (oFFStop[85]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[85])
);

(* LOC = "SLICE_X87Y132" *)
      FDCE #(.INIT(1'b0)) Stopff86(
          .Q          (oFFStop[86]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[86])
);

(* LOC = "SLICE_X87Y132" *)
      FDCE #(.INIT(1'b0)) Stopff87(
          .Q          (oFFStop[87]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[87])
);

(* LOC = "SLICE_X87Y133" *)
      FDCE #(.INIT(1'b0)) Stopff88(
          .Q          (oFFStop[88]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[88])
);

(* LOC = "SLICE_X87Y133" *)
      FDCE #(.INIT(1'b0)) Stopff89(
          .Q          (oFFStop[89]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[89])
);

(* LOC = "SLICE_X87Y133" *)
      FDCE #(.INIT(1'b0)) Stopff90(
          .Q          (oFFStop[90]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[90])
);

(* LOC = "SLICE_X87Y133" *)
      FDCE #(.INIT(1'b0)) Stopff91(
          .Q          (oFFStop[91]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[91])
);

(* LOC = "SLICE_X87Y134" *)
      FDCE #(.INIT(1'b0)) Stopff92(
          .Q          (oFFStop[92]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[92])
);

(* LOC = "SLICE_X87Y134" *)
      FDCE #(.INIT(1'b0)) Stopff93(
          .Q          (oFFStop[93]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[93])
);

(* LOC = "SLICE_X87Y134" *)
      FDCE #(.INIT(1'b0)) Stopff94(
          .Q          (oFFStop[94]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[94])
);

(* LOC = "SLICE_X87Y134" *)
      FDCE #(.INIT(1'b0)) Stopff95(
          .Q          (oFFStop[95]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[95])
);

(* LOC = "SLICE_X87Y135" *)
      FDCE #(.INIT(1'b0)) Stopff96(
          .Q          (oFFStop[96]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[96])
);

(* LOC = "SLICE_X87Y135" *)
      FDCE #(.INIT(1'b0)) Stopff97(
          .Q          (oFFStop[97]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[97])
);

(* LOC = "SLICE_X87Y135" *)
      FDCE #(.INIT(1'b0)) Stopff98(
          .Q          (oFFStop[98]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[98])
);

(* LOC = "SLICE_X87Y135" *)
      FDCE #(.INIT(1'b0)) Stopff99(
          .Q          (oFFStop[99]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[99])
);

(* LOC = "SLICE_X87Y136" *)
      FDCE #(.INIT(1'b0)) Stopff100(
          .Q          (oFFStop[100]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[100])
);

(* LOC = "SLICE_X87Y136" *)
      FDCE #(.INIT(1'b0)) Stopff101(
          .Q          (oFFStop[101]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[101])
);

(* LOC = "SLICE_X87Y136" *)
      FDCE #(.INIT(1'b0)) Stopff102(
          .Q          (oFFStop[102]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[102])
);

(* LOC = "SLICE_X87Y136" *)
      FDCE #(.INIT(1'b0)) Stopff103(
          .Q          (oFFStop[103]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[103])
);

(* LOC = "SLICE_X87Y137" *)
      FDCE #(.INIT(1'b0)) Stopff104(
          .Q          (oFFStop[104]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[104])
);

(* LOC = "SLICE_X87Y137" *)
      FDCE #(.INIT(1'b0)) Stopff105(
          .Q          (oFFStop[105]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[105])
);

(* LOC = "SLICE_X87Y137" *)
      FDCE #(.INIT(1'b0)) Stopff106(
          .Q          (oFFStop[106]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[106])
);

(* LOC = "SLICE_X87Y137" *)
      FDCE #(.INIT(1'b0)) Stopff107(
          .Q          (oFFStop[107]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[107])
);

(* LOC = "SLICE_X87Y138" *)
      FDCE #(.INIT(1'b0)) Stopff108(
          .Q          (oFFStop[108]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[108])
);

(* LOC = "SLICE_X87Y138" *)
      FDCE #(.INIT(1'b0)) Stopff109(
          .Q          (oFFStop[109]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[109])
);

(* LOC = "SLICE_X87Y138" *)
      FDCE #(.INIT(1'b0)) Stopff110(
          .Q          (oFFStop[110]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[110])
);

(* LOC = "SLICE_X87Y138" *)
      FDCE #(.INIT(1'b0)) Stopff111(
          .Q          (oFFStop[111]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[111])
);

(* LOC = "SLICE_X87Y139" *)
      FDCE #(.INIT(1'b0)) Stopff112(
          .Q          (oFFStop[112]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[112])
);

(* LOC = "SLICE_X87Y139" *)
      FDCE #(.INIT(1'b0)) Stopff113(
          .Q          (oFFStop[113]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[113])
);

(* LOC = "SLICE_X87Y139" *)
      FDCE #(.INIT(1'b0)) Stopff114(
          .Q          (oFFStop[114]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[114])
);

(* LOC = "SLICE_X87Y139" *)
      FDCE #(.INIT(1'b0)) Stopff115(
          .Q          (oFFStop[115]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[115])
);

(* LOC = "SLICE_X87Y140" *)
      FDCE #(.INIT(1'b0)) Stopff116(
          .Q          (oFFStop[116]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[116])
);

(* LOC = "SLICE_X87Y140" *)
      FDCE #(.INIT(1'b0)) Stopff117(
          .Q          (oFFStop[117]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[117])
);

(* LOC = "SLICE_X87Y140" *)
      FDCE #(.INIT(1'b0)) Stopff118(
          .Q          (oFFStop[118]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[118])
);

(* LOC = "SLICE_X87Y140" *)
      FDCE #(.INIT(1'b0)) Stopff119(
          .Q          (oFFStop[119]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[119])
);

(* LOC = "SLICE_X87Y141" *)
      FDCE #(.INIT(1'b0)) Stopff120(
          .Q          (oFFStop[120]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[120])
);

(* LOC = "SLICE_X87Y141" *)
      FDCE #(.INIT(1'b0)) Stopff121(
          .Q          (oFFStop[121]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[121])
);

(* LOC = "SLICE_X87Y141" *)
      FDCE #(.INIT(1'b0)) Stopff122(
          .Q          (oFFStop[122]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[122])
);

(* LOC = "SLICE_X87Y141" *)
      FDCE #(.INIT(1'b0)) Stopff123(
          .Q          (oFFStop[123]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[123])
);

(* LOC = "SLICE_X87Y142" *)
      FDCE #(.INIT(1'b0)) Stopff124(
          .Q          (oFFStop[124]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[124])
);

(* LOC = "SLICE_X87Y142" *)
      FDCE #(.INIT(1'b0)) Stopff125(
          .Q          (oFFStop[125]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[125])
);

(* LOC = "SLICE_X87Y142" *)
      FDCE #(.INIT(1'b0)) Stopff126(
          .Q          (oFFStop[126]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[126])
);

(* LOC = "SLICE_X87Y142" *)
      FDCE #(.INIT(1'b0)) Stopff127(
          .Q          (oFFStop[127]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[127])
);

(* LOC = "SLICE_X87Y143" *)
      FDCE #(.INIT(1'b0)) Stopff128(
          .Q          (oFFStop[128]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[128])
);

(* LOC = "SLICE_X87Y143" *)
      FDCE #(.INIT(1'b0)) Stopff129(
          .Q          (oFFStop[129]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[129])
);

(* LOC = "SLICE_X87Y143" *)
      FDCE #(.INIT(1'b0)) Stopff130(
          .Q          (oFFStop[130]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[130])
);

(* LOC = "SLICE_X87Y143" *)
      FDCE #(.INIT(1'b0)) Stopff131(
          .Q          (oFFStop[131]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[131])
);

(* LOC = "SLICE_X87Y144" *)
      FDCE #(.INIT(1'b0)) Stopff132(
          .Q          (oFFStop[132]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[132])
);

(* LOC = "SLICE_X87Y144" *)
      FDCE #(.INIT(1'b0)) Stopff133(
          .Q          (oFFStop[133]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[133])
);

(* LOC = "SLICE_X87Y144" *)
      FDCE #(.INIT(1'b0)) Stopff134(
          .Q          (oFFStop[134]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[134])
);

(* LOC = "SLICE_X87Y144" *)
      FDCE #(.INIT(1'b0)) Stopff135(
          .Q          (oFFStop[135]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[135])
);

(* LOC = "SLICE_X87Y145" *)
      FDCE #(.INIT(1'b0)) Stopff136(
          .Q          (oFFStop[136]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[136])
);

(* LOC = "SLICE_X87Y145" *)
      FDCE #(.INIT(1'b0)) Stopff137(
          .Q          (oFFStop[137]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[137])
);

(* LOC = "SLICE_X87Y145" *)
      FDCE #(.INIT(1'b0)) Stopff138(
          .Q          (oFFStop[138]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[138])
);

(* LOC = "SLICE_X87Y145" *)
      FDCE #(.INIT(1'b0)) Stopff139(
          .Q          (oFFStop[139]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[139])
);

(* LOC = "SLICE_X87Y146" *)
      FDCE #(.INIT(1'b0)) Stopff140(
          .Q          (oFFStop[140]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[140])
);

(* LOC = "SLICE_X87Y146" *)
      FDCE #(.INIT(1'b0)) Stopff141(
          .Q          (oFFStop[141]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[141])
);

(* LOC = "SLICE_X87Y146" *)
      FDCE #(.INIT(1'b0)) Stopff142(
          .Q          (oFFStop[142]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[142])
);

(* LOC = "SLICE_X87Y146" *)
      FDCE #(.INIT(1'b0)) Stopff143(
          .Q          (oFFStop[143]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[143])
);

(* LOC = "SLICE_X87Y147" *)
      FDCE #(.INIT(1'b0)) Stopff144(
          .Q          (oFFStop[144]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[144])
);

(* LOC = "SLICE_X87Y147" *)
      FDCE #(.INIT(1'b0)) Stopff145(
          .Q          (oFFStop[145]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[145])
);

(* LOC = "SLICE_X87Y147" *)
      FDCE #(.INIT(1'b0)) Stopff146(
          .Q          (oFFStop[146]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[146])
);

(* LOC = "SLICE_X87Y147" *)
      FDCE #(.INIT(1'b0)) Stopff147(
          .Q          (oFFStop[147]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[147])
);

(* LOC = "SLICE_X87Y148" *)
      FDCE #(.INIT(1'b0)) Stopff148(
          .Q          (oFFStop[148]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[148])
);

(* LOC = "SLICE_X87Y148" *)
      FDCE #(.INIT(1'b0)) Stopff149(
          .Q          (oFFStop[149]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[149])
);

(* LOC = "SLICE_X87Y148" *)
      FDCE #(.INIT(1'b0)) Stopff150(
          .Q          (oFFStop[150]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[150])
);

(* LOC = "SLICE_X87Y148" *)
      FDCE #(.INIT(1'b0)) Stopff151(
          .Q          (oFFStop[151]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[151])
);

(* LOC = "SLICE_X87Y149" *)
      FDCE #(.INIT(1'b0)) Stopff152(
          .Q          (oFFStop[152]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[152])
);

(* LOC = "SLICE_X87Y149" *)
      FDCE #(.INIT(1'b0)) Stopff153(
          .Q          (oFFStop[153]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[153])
);

(* LOC = "SLICE_X87Y149" *)
      FDCE #(.INIT(1'b0)) Stopff154(
          .Q          (oFFStop[154]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[154])
);

(* LOC = "SLICE_X87Y149" *)
      FDCE #(.INIT(1'b0)) Stopff155(
          .Q          (oFFStop[155]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[155])
);

(* LOC = "SLICE_X87Y150" *)
      FDCE #(.INIT(1'b0)) Stopff156(
          .Q          (oFFStop[156]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[156])
);

(* LOC = "SLICE_X87Y150" *)
      FDCE #(.INIT(1'b0)) Stopff157(
          .Q          (oFFStop[157]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[157])
);

(* LOC = "SLICE_X87Y150" *)
      FDCE #(.INIT(1'b0)) Stopff158(
          .Q          (oFFStop[158]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[158])
);

(* LOC = "SLICE_X87Y150" *)
      FDCE #(.INIT(1'b0)) Stopff159(
          .Q          (oFFStop[159]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[159])
);

(* LOC = "SLICE_X87Y151" *)
      FDCE #(.INIT(1'b0)) Stopff160(
          .Q          (oFFStop[160]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[160])
);

(* LOC = "SLICE_X87Y151" *)
      FDCE #(.INIT(1'b0)) Stopff161(
          .Q          (oFFStop[161]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[161])
);

(* LOC = "SLICE_X87Y151" *)
      FDCE #(.INIT(1'b0)) Stopff162(
          .Q          (oFFStop[162]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[162])
);

(* LOC = "SLICE_X87Y151" *)
      FDCE #(.INIT(1'b0)) Stopff163(
          .Q          (oFFStop[163]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[163])
);

(* LOC = "SLICE_X87Y152" *)
      FDCE #(.INIT(1'b0)) Stopff164(
          .Q          (oFFStop[164]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[164])
);

(* LOC = "SLICE_X87Y152" *)
      FDCE #(.INIT(1'b0)) Stopff165(
          .Q          (oFFStop[165]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[165])
);

(* LOC = "SLICE_X87Y152" *)
      FDCE #(.INIT(1'b0)) Stopff166(
          .Q          (oFFStop[166]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[166])
);

(* LOC = "SLICE_X87Y152" *)
      FDCE #(.INIT(1'b0)) Stopff167(
          .Q          (oFFStop[167]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[167])
);

(* LOC = "SLICE_X87Y153" *)
      FDCE #(.INIT(1'b0)) Stopff168(
          .Q          (oFFStop[168]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[168])
);

(* LOC = "SLICE_X87Y153" *)
      FDCE #(.INIT(1'b0)) Stopff169(
          .Q          (oFFStop[169]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[169])
);

(* LOC = "SLICE_X87Y153" *)
      FDCE #(.INIT(1'b0)) Stopff170(
          .Q          (oFFStop[170]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[170])
);

(* LOC = "SLICE_X87Y153" *)
      FDCE #(.INIT(1'b0)) Stopff171(
          .Q          (oFFStop[171]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[171])
);

(* LOC = "SLICE_X87Y154" *)
      FDCE #(.INIT(1'b0)) Stopff172(
          .Q          (oFFStop[172]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[172])
);

(* LOC = "SLICE_X87Y154" *)
      FDCE #(.INIT(1'b0)) Stopff173(
          .Q          (oFFStop[173]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[173])
);

(* LOC = "SLICE_X87Y154" *)
      FDCE #(.INIT(1'b0)) Stopff174(
          .Q          (oFFStop[174]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[174])
);

(* LOC = "SLICE_X87Y154" *)
      FDCE #(.INIT(1'b0)) Stopff175(
          .Q          (oFFStop[175]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[175])
);

(* LOC = "SLICE_X87Y155" *)
      FDCE #(.INIT(1'b0)) Stopff176(
          .Q          (oFFStop[176]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[176])
);

(* LOC = "SLICE_X87Y155" *)
      FDCE #(.INIT(1'b0)) Stopff177(
          .Q          (oFFStop[177]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[177])
);

(* LOC = "SLICE_X87Y155" *)
      FDCE #(.INIT(1'b0)) Stopff178(
          .Q          (oFFStop[178]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[178])
);

(* LOC = "SLICE_X87Y155" *)
      FDCE #(.INIT(1'b0)) Stopff179(
          .Q          (oFFStop[179]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[179])
);

(* LOC = "SLICE_X87Y156" *)
      FDCE #(.INIT(1'b0)) Stopff180(
          .Q          (oFFStop[180]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[180])
);

(* LOC = "SLICE_X87Y156" *)
      FDCE #(.INIT(1'b0)) Stopff181(
          .Q          (oFFStop[181]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[181])
);

(* LOC = "SLICE_X87Y156" *)
      FDCE #(.INIT(1'b0)) Stopff182(
          .Q          (oFFStop[182]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[182])
);

(* LOC = "SLICE_X87Y156" *)
      FDCE #(.INIT(1'b0)) Stopff183(
          .Q          (oFFStop[183]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[183])
);

(* LOC = "SLICE_X87Y157" *)
      FDCE #(.INIT(1'b0)) Stopff184(
          .Q          (oFFStop[184]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[184])
);

(* LOC = "SLICE_X87Y157" *)
      FDCE #(.INIT(1'b0)) Stopff185(
          .Q          (oFFStop[185]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[185])
);

(* LOC = "SLICE_X87Y157" *)
      FDCE #(.INIT(1'b0)) Stopff186(
          .Q          (oFFStop[186]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[186])
);

(* LOC = "SLICE_X87Y157" *)
      FDCE #(.INIT(1'b0)) Stopff187(
          .Q          (oFFStop[187]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[187])
);

(* LOC = "SLICE_X87Y158" *)
      FDCE #(.INIT(1'b0)) Stopff188(
          .Q          (oFFStop[188]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[188])
);

(* LOC = "SLICE_X87Y158" *)
      FDCE #(.INIT(1'b0)) Stopff189(
          .Q          (oFFStop[189]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[189])
);

(* LOC = "SLICE_X87Y158" *)
      FDCE #(.INIT(1'b0)) Stopff190(
          .Q          (oFFStop[190]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[190])
);

(* LOC = "SLICE_X87Y158" *)
      FDCE #(.INIT(1'b0)) Stopff191(
          .Q          (oFFStop[191]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[191])
);

(* LOC = "SLICE_X87Y159" *)
      FDCE #(.INIT(1'b0)) Stopff192(
          .Q          (oFFStop[192]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[192])
);

(* LOC = "SLICE_X87Y159" *)
      FDCE #(.INIT(1'b0)) Stopff193(
          .Q          (oFFStop[193]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[193])
);

(* LOC = "SLICE_X87Y159" *)
      FDCE #(.INIT(1'b0)) Stopff194(
          .Q          (oFFStop[194]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[194])
);

(* LOC = "SLICE_X87Y159" *)
      FDCE #(.INIT(1'b0)) Stopff195(
          .Q          (oFFStop[195]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[195])
);

(* LOC = "SLICE_X87Y160" *)
      FDCE #(.INIT(1'b0)) Stopff196(
          .Q          (oFFStop[196]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[196])
);

(* LOC = "SLICE_X87Y160" *)
      FDCE #(.INIT(1'b0)) Stopff197(
          .Q          (oFFStop[197]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[197])
);

(* LOC = "SLICE_X87Y160" *)
      FDCE #(.INIT(1'b0)) Stopff198(
          .Q          (oFFStop[198]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[198])
);

(* LOC = "SLICE_X87Y160" *)
      FDCE #(.INIT(1'b0)) Stopff199(
          .Q          (oFFStop[199]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[199])
);

(* LOC = "SLICE_X87Y161" *)
      FDCE #(.INIT(1'b0)) Stopff200(
          .Q          (oFFStop[200]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[200])
);

(* LOC = "SLICE_X87Y161" *)
      FDCE #(.INIT(1'b0)) Stopff201(
          .Q          (oFFStop[201]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[201])
);

(* LOC = "SLICE_X87Y161" *)
      FDCE #(.INIT(1'b0)) Stopff202(
          .Q          (oFFStop[202]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[202])
);

(* LOC = "SLICE_X87Y161" *)
      FDCE #(.INIT(1'b0)) Stopff203(
          .Q          (oFFStop[203]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[203])
);

(* LOC = "SLICE_X87Y162" *)
      FDCE #(.INIT(1'b0)) Stopff204(
          .Q          (oFFStop[204]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[204])
);

(* LOC = "SLICE_X87Y162" *)
      FDCE #(.INIT(1'b0)) Stopff205(
          .Q          (oFFStop[205]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[205])
);

(* LOC = "SLICE_X87Y162" *)
      FDCE #(.INIT(1'b0)) Stopff206(
          .Q          (oFFStop[206]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[206])
);

(* LOC = "SLICE_X87Y162" *)
      FDCE #(.INIT(1'b0)) Stopff207(
          .Q          (oFFStop[207]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[207])
);

(* LOC = "SLICE_X87Y163" *)
      FDCE #(.INIT(1'b0)) Stopff208(
          .Q          (oFFStop[208]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[208])
);

(* LOC = "SLICE_X87Y163" *)
      FDCE #(.INIT(1'b0)) Stopff209(
          .Q          (oFFStop[209]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[209])
);

(* LOC = "SLICE_X87Y163" *)
      FDCE #(.INIT(1'b0)) Stopff210(
          .Q          (oFFStop[210]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[210])
);

(* LOC = "SLICE_X87Y163" *)
      FDCE #(.INIT(1'b0)) Stopff211(
          .Q          (oFFStop[211]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[211])
);

(* LOC = "SLICE_X87Y164" *)
      FDCE #(.INIT(1'b0)) Stopff212(
          .Q          (oFFStop[212]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[212])
);

(* LOC = "SLICE_X87Y164" *)
      FDCE #(.INIT(1'b0)) Stopff213(
          .Q          (oFFStop[213]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[213])
);

(* LOC = "SLICE_X87Y164" *)
      FDCE #(.INIT(1'b0)) Stopff214(
          .Q          (oFFStop[214]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[214])
);

(* LOC = "SLICE_X87Y164" *)
      FDCE #(.INIT(1'b0)) Stopff215(
          .Q          (oFFStop[215]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[215])
);

(* LOC = "SLICE_X87Y165" *)
      FDCE #(.INIT(1'b0)) Stopff216(
          .Q          (oFFStop[216]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[216])
);

(* LOC = "SLICE_X87Y165" *)
      FDCE #(.INIT(1'b0)) Stopff217(
          .Q          (oFFStop[217]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[217])
);

(* LOC = "SLICE_X87Y165" *)
      FDCE #(.INIT(1'b0)) Stopff218(
          .Q          (oFFStop[218]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[218])
);

(* LOC = "SLICE_X87Y165" *)
      FDCE #(.INIT(1'b0)) Stopff219(
          .Q          (oFFStop[219]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[219])
);

(* LOC = "SLICE_X87Y166" *)
      FDCE #(.INIT(1'b0)) Stopff220(
          .Q          (oFFStop[220]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[220])
);

(* LOC = "SLICE_X87Y166" *)
      FDCE #(.INIT(1'b0)) Stopff221(
          .Q          (oFFStop[221]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[221])
);

(* LOC = "SLICE_X87Y166" *)
      FDCE #(.INIT(1'b0)) Stopff222(
          .Q          (oFFStop[222]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[222])
);

(* LOC = "SLICE_X87Y166" *)
      FDCE #(.INIT(1'b0)) Stopff223(
          .Q          (oFFStop[223]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[223])
);

(* LOC = "SLICE_X87Y167" *)
      FDCE #(.INIT(1'b0)) Stopff224(
          .Q          (oFFStop[224]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[224])
);

(* LOC = "SLICE_X87Y167" *)
      FDCE #(.INIT(1'b0)) Stopff225(
          .Q          (oFFStop[225]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[225])
);

(* LOC = "SLICE_X87Y167" *)
      FDCE #(.INIT(1'b0)) Stopff226(
          .Q          (oFFStop[226]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[226])
);

(* LOC = "SLICE_X87Y167" *)
      FDCE #(.INIT(1'b0)) Stopff227(
          .Q          (oFFStop[227]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[227])
);

(* LOC = "SLICE_X87Y168" *)
      FDCE #(.INIT(1'b0)) Stopff228(
          .Q          (oFFStop[228]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[228])
);

(* LOC = "SLICE_X87Y168" *)
      FDCE #(.INIT(1'b0)) Stopff229(
          .Q          (oFFStop[229]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[229])
);

(* LOC = "SLICE_X87Y168" *)
      FDCE #(.INIT(1'b0)) Stopff230(
          .Q          (oFFStop[230]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[230])
);

(* LOC = "SLICE_X87Y168" *)
      FDCE #(.INIT(1'b0)) Stopff231(
          .Q          (oFFStop[231]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[231])
);

(* LOC = "SLICE_X87Y169" *)
      FDCE #(.INIT(1'b0)) Stopff232(
          .Q          (oFFStop[232]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[232])
);

(* LOC = "SLICE_X87Y169" *)
      FDCE #(.INIT(1'b0)) Stopff233(
          .Q          (oFFStop[233]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[233])
);

(* LOC = "SLICE_X87Y169" *)
      FDCE #(.INIT(1'b0)) Stopff234(
          .Q          (oFFStop[234]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[234])
);

(* LOC = "SLICE_X87Y169" *)
      FDCE #(.INIT(1'b0)) Stopff235(
          .Q          (oFFStop[235]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[235])
);

(* LOC = "SLICE_X87Y170" *)
      FDCE #(.INIT(1'b0)) Stopff236(
          .Q          (oFFStop[236]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[236])
);

(* LOC = "SLICE_X87Y170" *)
      FDCE #(.INIT(1'b0)) Stopff237(
          .Q          (oFFStop[237]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[237])
);

(* LOC = "SLICE_X87Y170" *)
      FDCE #(.INIT(1'b0)) Stopff238(
          .Q          (oFFStop[238]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[238])
);

(* LOC = "SLICE_X87Y170" *)
      FDCE #(.INIT(1'b0)) Stopff239(
          .Q          (oFFStop[239]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[239])
);

(* LOC = "SLICE_X87Y171" *)
      FDCE #(.INIT(1'b0)) Stopff240(
          .Q          (oFFStop[240]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[240])
);

(* LOC = "SLICE_X87Y171" *)
      FDCE #(.INIT(1'b0)) Stopff241(
          .Q          (oFFStop[241]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[241])
);

(* LOC = "SLICE_X87Y171" *)
      FDCE #(.INIT(1'b0)) Stopff242(
          .Q          (oFFStop[242]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[242])
);

(* LOC = "SLICE_X87Y171" *)
      FDCE #(.INIT(1'b0)) Stopff243(
          .Q          (oFFStop[243]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[243])
);

(* LOC = "SLICE_X87Y172" *)
      FDCE #(.INIT(1'b0)) Stopff244(
          .Q          (oFFStop[244]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[244])
);

(* LOC = "SLICE_X87Y172" *)
      FDCE #(.INIT(1'b0)) Stopff245(
          .Q          (oFFStop[245]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[245])
);

(* LOC = "SLICE_X87Y172" *)
      FDCE #(.INIT(1'b0)) Stopff246(
          .Q          (oFFStop[246]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[246])
);

(* LOC = "SLICE_X87Y172" *)
      FDCE #(.INIT(1'b0)) Stopff247(
          .Q          (oFFStop[247]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[247])
);

(* LOC = "SLICE_X87Y173" *)
      FDCE #(.INIT(1'b0)) Stopff248(
          .Q          (oFFStop[248]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[248])
);

(* LOC = "SLICE_X87Y173" *)
      FDCE #(.INIT(1'b0)) Stopff249(
          .Q          (oFFStop[249]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[249])
);

(* LOC = "SLICE_X87Y173" *)
      FDCE #(.INIT(1'b0)) Stopff250(
          .Q          (oFFStop[250]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[250])
);

(* LOC = "SLICE_X87Y173" *)
      FDCE #(.INIT(1'b0)) Stopff251(
          .Q          (oFFStop[251]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[251])
);

(* LOC = "SLICE_X87Y174" *)
      FDCE #(.INIT(1'b0)) Stopff252(
          .Q          (oFFStop[252]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[252])
);

(* LOC = "SLICE_X87Y174" *)
      FDCE #(.INIT(1'b0)) Stopff253(
          .Q          (oFFStop[253]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[253])
);

(* LOC = "SLICE_X87Y174" *)
      FDCE #(.INIT(1'b0)) Stopff254(
          .Q          (oFFStop[254]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[254])
);

(* LOC = "SLICE_X87Y174" *)
      FDCE #(.INIT(1'b0)) Stopff255(
          .Q          (oFFStop[255]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[255])
);

(* LOC = "SLICE_X87Y175" *)
      FDCE #(.INIT(1'b0)) Stopff256(
          .Q          (oFFStop[256]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[256])
);

(* LOC = "SLICE_X87Y175" *)
      FDCE #(.INIT(1'b0)) Stopff257(
          .Q          (oFFStop[257]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[257])
);

(* LOC = "SLICE_X87Y175" *)
      FDCE #(.INIT(1'b0)) Stopff258(
          .Q          (oFFStop[258]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[258])
);

(* LOC = "SLICE_X87Y175" *)
      FDCE #(.INIT(1'b0)) Stopff259(
          .Q          (oFFStop[259]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[259])
);

(* LOC = "SLICE_X87Y176" *)
      FDCE #(.INIT(1'b0)) Stopff260(
          .Q          (oFFStop[260]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[260])
);

(* LOC = "SLICE_X87Y176" *)
      FDCE #(.INIT(1'b0)) Stopff261(
          .Q          (oFFStop[261]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[261])
);

(* LOC = "SLICE_X87Y176" *)
      FDCE #(.INIT(1'b0)) Stopff262(
          .Q          (oFFStop[262]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[262])
);

(* LOC = "SLICE_X87Y176" *)
      FDCE #(.INIT(1'b0)) Stopff263(
          .Q          (oFFStop[263]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[263])
);

(* LOC = "SLICE_X87Y177" *)
      FDCE #(.INIT(1'b0)) Stopff264(
          .Q          (oFFStop[264]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[264])
);

(* LOC = "SLICE_X87Y177" *)
      FDCE #(.INIT(1'b0)) Stopff265(
          .Q          (oFFStop[265]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[265])
);

(* LOC = "SLICE_X87Y177" *)
      FDCE #(.INIT(1'b0)) Stopff266(
          .Q          (oFFStop[266]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[266])
);

(* LOC = "SLICE_X87Y177" *)
      FDCE #(.INIT(1'b0)) Stopff267(
          .Q          (oFFStop[267]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[267])
);

(* LOC = "SLICE_X87Y178" *)
      FDCE #(.INIT(1'b0)) Stopff268(
          .Q          (oFFStop[268]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[268])
);

(* LOC = "SLICE_X87Y178" *)
      FDCE #(.INIT(1'b0)) Stopff269(
          .Q          (oFFStop[269]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[269])
);

(* LOC = "SLICE_X87Y178" *)
      FDCE #(.INIT(1'b0)) Stopff270(
          .Q          (oFFStop[270]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[270])
);

(* LOC = "SLICE_X87Y178" *)
      FDCE #(.INIT(1'b0)) Stopff271(
          .Q          (oFFStop[271]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[271])
);

(* LOC = "SLICE_X87Y179" *)
      FDCE #(.INIT(1'b0)) Stopff272(
          .Q          (oFFStop[272]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[272])
);

(* LOC = "SLICE_X87Y179" *)
      FDCE #(.INIT(1'b0)) Stopff273(
          .Q          (oFFStop[273]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[273])
);

(* LOC = "SLICE_X87Y179" *)
      FDCE #(.INIT(1'b0)) Stopff274(
          .Q          (oFFStop[274]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[274])
);

(* LOC = "SLICE_X87Y179" *)
      FDCE #(.INIT(1'b0)) Stopff275(
          .Q          (oFFStop[275]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[275])
);

(* LOC = "SLICE_X87Y180" *)
      FDCE #(.INIT(1'b0)) Stopff276(
          .Q          (oFFStop[276]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[276])
);

(* LOC = "SLICE_X87Y180" *)
      FDCE #(.INIT(1'b0)) Stopff277(
          .Q          (oFFStop[277]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[277])
);

(* LOC = "SLICE_X87Y180" *)
      FDCE #(.INIT(1'b0)) Stopff278(
          .Q          (oFFStop[278]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[278])
);

(* LOC = "SLICE_X87Y180" *)
      FDCE #(.INIT(1'b0)) Stopff279(
          .Q          (oFFStop[279]),
          .C          (clk),
          .CE         (iStopEnable),
          .CLR        (iRst),
          .D          (wFirstFF[279])
);

endmodule //
