//////////////////////////////////////////////////////////////////////
// Module Name: decode_tb
// 
//
// Author: Miqueas Filsinger
// Date: 03-06-2024
//
// Revision History:
// 
// Notes:
// - Any additional notes or considerations
//
//////////////////////////////////////////////////////////////////////

module decode_tb (
    // Ports here
);

    

endmodule //