//////////////////////////////////////////////////////////////////////
// Module Name: Decoder
// Description: Brief description of the module's functionality
//
// Author: Miqueas Filsinger
// Date: Date Created or Last Modified
//
// Revision History:
// - Date: Description of changes made
// - Date: Description of changes made
//
// Notes:
// - Any additional notes or considerations
//
//////////////////////////////////////////////////////////////////////

module Decoder #(parameter NUM = 12)(
    input  wire[NUM-1:0]    iFF
);

    
endmodule //