//////////////////////////////////////////////////////////////////////
// Module Name: Input
// Description: Settle Wave Union A (WU-A) principles to source the Fine delay chain.
//
// Author: Miqueas Filsinger
// Date: Date 
//
// Revision History:
//
// Notes:
// - 
//
//////////////////////////////////////////////////////////////////////

module  Input(
    // Ports here
);

    // Module implementation here

endmodule //